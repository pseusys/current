�� sr java.util.HashMap���`� F 
loadFactorI 	thresholdxp?@     w      t NODESsq ~  ?@     w      
sr java.lang.Integer⠤���8 I valuexr java.lang.Number������  xp    sq ~  ?@     w      t POSITIONsr java.lang.Boolean� r�՜�� Z valuexpt ARKSsq ~  ?@     w      q ~ sq ~  ?@     w      t STARTt At ENDt Lt HIDDENq ~ 
t WEIGHTsr java.lang.Double���J)k� D valuexq ~ @       xsq ~    sq ~  ?@     w      q ~ q ~ q ~ t Gq ~ q ~ 
q ~ sq ~ @      xsq ~    sq ~  ?@     w      q ~ q ~ q ~ t Hq ~ q ~ 
q ~ sq ~ @      xxt 
POSITION_Xsq ~ @s`     t 
POSITION_Ysq ~ @s�     q ~ q ~ 
t NAMEq ~ xq ~ sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ t Dq ~ q ~ q ~ q ~ 
q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ q ~ t Fq ~ q ~ 
q ~ sq ~ @      xxq ~ sq ~ @�     q ~  sq ~ @|0     q ~ q ~ 
q ~ "q ~ xq ~ sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ t Cq ~ q ~ q ~ q ~ 
q ~ sq ~ @7      xq ~ sq ~  ?@     w      q ~ q ~ q ~ t Qq ~ q ~ 
q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ @      xxq ~ sq ~ @�      q ~  sq ~ @s�     q ~ q ~ 
q ~ "q ~ xsq ~    sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ t Bq ~ q ~ +q ~ q ~ 
q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ 5q ~ q ~ +q ~ q ~ 
q ~ sq ~ @       xq ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ +q ~ q ~ 
q ~ sq ~ @      xxq ~ sq ~ @z�     q ~  sq ~ @k@     q ~ q ~ 
q ~ "q ~ +xsq ~    sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ q ~ t Eq ~ q ~ 
q ~ sq ~ @&      xq ~ sq ~  ?@     w      q ~ q ~ 5q ~ q ~ Kq ~ q ~ 
q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ &q ~ q ~ Kq ~ q ~ 
q ~ sq ~ @4      xxq ~ sq ~ @p     q ~  sq ~ @��     q ~ q ~ 
q ~ "q ~ Kxsq ~    sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ &q ~ q ~ 2q ~ q ~ 
q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ &q ~ q ~ Kq ~ q ~ 
q ~ sq ~ @4      xq ~ sq ~  ?@     w      q ~ q ~ &q ~ q ~ q ~ q ~ 
q ~ sq ~ @      xxq ~ sq ~ @�h     q ~  sq ~ @��     q ~ q ~ 
q ~ "q ~ &xsq ~    sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ 2q ~ q ~ ?q ~ q ~ 
q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ 2q ~ q ~ q ~ q ~ 
q ~ sq ~ @7      xq ~ sq ~  ?@     w      q ~ q ~ &q ~ q ~ 2q ~ q ~ 
q ~ sq ~ @      xxq ~ sq ~ @��     q ~  sq ~ @r�     q ~ q ~ 
q ~ "q ~ 2xsq ~    sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ ?q ~ q ~ q ~ q ~ 
q ~ sq ~ @$      xq ~ sq ~  ?@     w      q ~ q ~ ?q ~ q ~ +q ~ q ~ 
q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ 2q ~ q ~ ?q ~ q ~ 
q ~ sq ~ @      xxq ~ sq ~ @{      q ~  sq ~ @T�     q ~ q ~ 
q ~ "q ~ ?xsq ~    sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ 5q ~ q ~ Kq ~ q ~ 
q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ 5q ~ q ~ +q ~ q ~ 
q ~ sq ~ @       xq ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ 5q ~ q ~ 
q ~ sq ~ @      xxq ~ sq ~ @u�     q ~  sq ~ @|@     q ~ q ~ 
q ~ "q ~ 5xsq ~    	sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ ?q ~ q ~ q ~ q ~ 
q ~ sq ~ @$      xq ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ Kq ~ q ~ 
q ~ sq ~ @&      xq ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ @       xxq ~ sq ~ @e�     q ~  sq ~ @r`     q ~ q ~ 
q ~ "q ~ xxq ~ sq ~  ?@     w       q ~ sq ~  ?@     w      q ~ q ~ ?q ~ q ~ q ~ q ~ 
q ~ sq ~ @$      xq ~ sq ~  ?@     w      q ~ q ~ ?q ~ q ~ +q ~ q ~ 
q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ 2q ~ q ~ ?q ~ q ~ 
q ~ sq ~ @      xq ~ ;sq ~  ?@     w      q ~ q ~ 2q ~ q ~ q ~ q ~ 
q ~ sq ~ @7      xq ~ Gsq ~  ?@     w      q ~ q ~ q ~ q ~ Kq ~ q ~ 
q ~ sq ~ @&      xq ~ Ssq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ @       xq ~ ^sq ~  ?@     w      q ~ q ~ 5q ~ q ~ Kq ~ q ~ 
q ~ sq ~ @      xq ~ isq ~  ?@     w      q ~ q ~ &q ~ q ~ 2q ~ q ~ 
q ~ sq ~ @      xq ~ tsq ~  ?@     w      q ~ q ~ &q ~ q ~ Kq ~ q ~ 
q ~ sq ~ @4      xq ~ sq ~  ?@     w      q ~ q ~ &q ~ q ~ q ~ q ~ 
q ~ sq ~ @      xsq ~    
sq ~  ?@     w      q ~ q ~ 5q ~ q ~ +q ~ q ~ 
q ~ sq ~ @       xsq ~    sq ~  ?@     w      q ~ q ~ q ~ q ~ 5q ~ q ~ 
q ~ sq ~ @      xsq ~    sq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ @      xsq ~    sq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ @      xsq ~    sq ~  ?@     w      q ~ q ~ q ~ q ~ +q ~ q ~ 
q ~ sq ~ @      xxx