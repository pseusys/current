�� sr java.util.HashMap���`� F 
loadFactorI 	thresholdxp?@     w      t NODESsq ~  ?@     w      sr java.lang.Integer⠤���8 I valuexr java.lang.Number������  xp    sq ~  ?@     w      t POSITIONsr java.lang.Boolean� r�՜�� Z valuexpt ARKSsq ~  ?@     w      q ~ sq ~  ?@     w      t STARTt Bt ENDt Gt HIDDENq ~ 
t WEIGHTsr java.lang.Double���J)k� D valuexq ~ @      xsq ~    sq ~  ?@     w      q ~ q ~ q ~ t Aq ~ sq ~ 	 q ~ sq ~ @       xsq ~    sq ~  ?@     w      q ~ t Cq ~ q ~ q ~ q ~ 
q ~ sq ~ @5      xxt 
POSITION_Xsq ~ @�P     t 
POSITION_Ysq ~ @��     q ~ q ~ 
t NAMEq ~ xq ~ sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ q ~ t Fq ~ q ~ q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ 'q ~ q ~ q ~ q ~ q ~ sq ~ @$      xxq ~ sq ~ @�(     q ~ !sq ~ @~�     q ~ q ~ 
q ~ #q ~ 'xq ~ sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ q ~ t Eq ~ q ~ q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ 0q ~ q ~ q ~ q ~ q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ 0q ~ q ~ 
q ~ sq ~ @$      xxq ~ sq ~ @��     q ~ !sq ~ @p`     q ~ q ~ 
q ~ #q ~ 0xsq ~    sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ q ~ t Dq ~ q ~ q ~ sq ~ @*      xxq ~ sq ~ @�8     q ~ !sq ~ @T@     q ~ q ~ 
q ~ #q ~ <xsq ~    sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ 'q ~ q ~ q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ @5      xq ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ 0q ~ q ~ 
q ~ sq ~ @$      xxq ~ sq ~ @e�     q ~ !sq ~ @��     q ~ q ~ 
q ~ #q ~ xsq ~    sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ 0q ~ q ~ q ~ q ~ q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ @      xxq ~ sq ~ @e�     q ~ !sq ~ @y      q ~ q ~ 
q ~ #q ~ xsq ~    sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ <q ~ q ~ q ~ sq ~ @*      xq ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ 0q ~ q ~ q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ q ~ sq ~ @       xq ~ 8sq ~  ?@     w      q ~ q ~ 'q ~ q ~ q ~ q ~ q ~ sq ~ @$      xxq ~ sq ~ @f      q ~ !sq ~ @n�     q ~ q ~ 
q ~ #q ~ xxq ~ sq ~  ?@     w      	q ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ <q ~ q ~ 
q ~ sq ~ @*      xq ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ 0q ~ q ~ 
q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ 0q ~ q ~ q ~ q ~ 
q ~ sq ~ @      xq ~ 8sq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ @      xq ~ @sq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ @       xq ~ Ksq ~  ?@     w      q ~ q ~ q ~ q ~ 'q ~ q ~ 
q ~ sq ~ @      xq ~ Tsq ~  ?@     w      q ~ q ~ 'q ~ q ~ q ~ q ~ 
q ~ sq ~ @$      xsq ~    sq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ @5      xsq ~    sq ~  ?@     w      q ~ q ~ q ~ q ~ 0q ~ q ~ 
q ~ sq ~ @$      xxx