�� sr java.util.HashMap���`� F 
loadFactorI 	thresholdxp?@     w      t NODESsq ~  ?@     w      sr java.lang.Integer⠤���8 I valuexr java.lang.Number������  xp    sq ~  ?@     w      t POSITIONsr java.lang.Boolean� r�՜�� Z valuexpt ARKSsq ~  ?@     w      q ~ sq ~  ?@     w      t STARTt At ENDt Ht HIDDENq ~ 
t WEIGHTsr java.lang.Double���J)k� D valuexq ~ @      xsq ~    sq ~  ?@     w      q ~ t Eq ~ q ~ q ~ q ~ 
q ~ sq ~ ?�      xxt 
POSITION_Xsq ~ @e�     t 
POSITION_Ysq ~ @u�     q ~ q ~ 
t NAMEq ~ xq ~ sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ q ~ t Gq ~ q ~ 
q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ t Fq ~ q ~ "q ~ q ~ 
q ~ sq ~ @       xxq ~ sq ~ @p�     q ~ sq ~ @�     q ~ q ~ 
q ~ q ~ "xsq ~    sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ %q ~ q ~ 
q ~ sq ~ @       xq ~ sq ~  ?@     w      q ~ q ~ %q ~ q ~ "q ~ q ~ 
q ~ sq ~ @       xq ~ )sq ~  ?@     w      q ~ t Dq ~ q ~ %q ~ q ~ 
q ~ sq ~ @      xxq ~ sq ~ @}@     q ~ sq ~ @��     q ~ q ~ 
q ~ q ~ %xsq ~    sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ ?�      xq ~ )sq ~  ?@     w      q ~ q ~ q ~ q ~ 1q ~ q ~ 
q ~ sq ~ @"      xxq ~ sq ~ @�     q ~ sq ~ @�p     q ~ q ~ 
q ~ q ~ xsq ~    sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ 1q ~ q ~ 
q ~ sq ~ @      xq ~ sq ~  ?@     w      q ~ q ~ 1q ~ t Bq ~ q ~ 
q ~ sq ~ @      xq ~ )sq ~  ?@     w      q ~ q ~ 1q ~ q ~ %q ~ q ~ 
q ~ sq ~ @      xq ~ 5sq ~  ?@     w      q ~ q ~ 1q ~ t Cq ~ q ~ 
q ~ sq ~ @*      xq ~ @sq ~  ?@     w      q ~ q ~ q ~ q ~ 1q ~ q ~ 
q ~ sq ~ @"      xxq ~ sq ~ @�X     q ~ sq ~ @vP     q ~ q ~ 
q ~ q ~ 1xsq ~    sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ Kq ~ q ~ 
q ~ sq ~ ?�      xq ~ sq ~  ?@     w      q ~ q ~ 1q ~ q ~ Kq ~ q ~ 
q ~ sq ~ @*      xxq ~ sq ~ @�h     q ~ sq ~ @g      q ~ q ~ 
q ~ q ~ Kxsq ~    sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ Fq ~ q ~ 
q ~ sq ~         xq ~ sq ~  ?@     w      q ~ q ~ 1q ~ q ~ Fq ~ q ~ 
q ~ sq ~ @      xxq ~ sq ~ @~`     q ~ sq ~ @]�     q ~ q ~ 
q ~ q ~ Fxsq ~    sq ~  ?@     w      q ~ q ~ 
q ~ sq ~  ?@     w      q ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ Fq ~ q ~ 
q ~ sq ~         xq ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ Kq ~ q ~ 
q ~ sq ~ ?�      xq ~ )sq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ @      xq ~ 5sq ~  ?@     w      q ~ q ~ q ~ q ~ 1q ~ q ~ 
q ~ sq ~ @      xq ~ @sq ~  ?@     w      q ~ q ~ q ~ q ~ %q ~ q ~ 
q ~ sq ~ @       xq ~ Qsq ~  ?@     w      q ~ q ~ q ~ q ~ "q ~ q ~ 
q ~ sq ~ @      xq ~ Zsq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ @      xxq ~ sq ~ @r�     q ~ sq ~ @e      q ~ q ~ 
q ~ q ~ xxq ~ sq ~  ?@     w       q ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ Fq ~ q ~ 
q ~ sq ~         xq ~ sq ~  ?@     w      q ~ q ~ q ~ q ~ Kq ~ q ~ 
q ~ sq ~ ?�      xq ~ )sq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ @      xq ~ 5sq ~  ?@     w      q ~ q ~ q ~ q ~ 1q ~ q ~ 
q ~ sq ~ @      xq ~ @sq ~  ?@     w      q ~ q ~ q ~ q ~ %q ~ q ~ 
q ~ sq ~ @       xq ~ Qsq ~  ?@     w      q ~ q ~ q ~ q ~ "q ~ q ~ 
q ~ sq ~ @      xq ~ Zsq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ @      xq ~ csq ~  ?@     w      q ~ q ~ %q ~ q ~ "q ~ q ~ 
q ~ sq ~ @       xsq ~    sq ~  ?@     w      q ~ q ~ 1q ~ q ~ Fq ~ q ~ 
q ~ sq ~ @      xsq ~    	sq ~  ?@     w      q ~ q ~ 1q ~ q ~ %q ~ q ~ 
q ~ sq ~ @      xsq ~    
sq ~  ?@     w      q ~ q ~ 1q ~ q ~ Kq ~ q ~ 
q ~ sq ~ @*      xsq ~    sq ~  ?@     w      q ~ q ~ q ~ q ~ q ~ q ~ 
q ~ sq ~ ?�      xsq ~    sq ~  ?@     w      q ~ q ~ q ~ q ~ 1q ~ q ~ 
q ~ sq ~ @"      xxx